/home/lunayang/Documents/Many-Core-SIMD-Research/lef/NangateOpenCellLibrary.lef