/home/lunayang/Documents/SIMAX/lef/NangateOpenCellLibrary.lef